// V, array length
// Tectonics: v run array-length.v
module main

// access array length
pub fn main() {
    arr := ["apple", "orange"]
    println(arr.len)
}
