module main;
  initial begin
    $display("0 ^ 0 = ", 0**0);
    $finish ;
  end
endmodule
