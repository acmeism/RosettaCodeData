module main;
  initial
    begin
      forever $display("SPAM");
    end
endmodule
