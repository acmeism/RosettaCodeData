import mymodule // name of module in those files

fn main() {
	mymodule.say_hi() // function from file 1 (myfile.v)
	mymodule.say_hi_and_bye() // function from file 2 (myfile2.v)
}
