// myfile.v
module mymodule

// Use "pub" to export a function
pub fn say_hi() {
	println("hello from mymodule!")
}
