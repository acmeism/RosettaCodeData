module main;
  initial begin
      $display("£");
    end
endmodule
