module mymodule

// To export a function we have to use `pub`

pub fn public_function() {
	println("hello from mymodule!")
}

fn private_function() {}
