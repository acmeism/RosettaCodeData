// Tokenize a string, in V (Vlang)
// Tectonics: v run tokenize-a-string.v
module main

// starts here
pub fn main() {
    println("Hello,How,Are,You,Today".split(',').join('.'))
}
