// Zero to the zero power, in V
// Tectonics: v run zero-to-the-zero-power.v
module main
import math

// starts here
// V does not include an exponentiation operator, but uses a math module
pub fn main() {
    println(math.pow(0, 0))
}
