module main;
  initial
    begin
      $write("Goodbye, World!");
      $finish ;
    end
endmodule
