module main
pub fn main() {}
