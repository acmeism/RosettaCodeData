entity dummy is
end;

architecture empty of dummy is
begin
end;
