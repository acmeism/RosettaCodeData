module mymodule

// To export a function we have to use 'pub'
pub fn say_hi() {
	println('hello from mymodule!')
}
