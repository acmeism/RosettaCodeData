module main;
endmodule
